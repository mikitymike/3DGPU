// $Id: $
// File name:   clip.sv
// Created:     4/29/2016
// Author:      Michael Malachowski
// Lab Section: 33704
// Version:     1.0  Initial Design Entry
// Description: Inputs a triangle, clips it, and outputs multiple triangles
