

module triangulizer
(
	input wire clk,
	input wire n_rst,
	input Polygon2D,


);

endmodule
