`ifndef CLIP_DEFINES_VH
`define CLIP_DEFINES_VH

`define INSIDE 'b0000
`define LEFT 'b0001
`define RIGHT 'b0010
`define BOTTOM 'b0100
`define TOP 'b1000
`define XMIN 0
`define XMAX 640
`define YMAX 480
`define YMIN 0

`endif